library verilog;
use verilog.vl_types.all;
entity clkgen_vlg_vec_tst is
end clkgen_vlg_vec_tst;
